`include "fifoCommon.sv"
`include "asyn_fifo.v"
`include "writeTx.sv"
`include "readTx.sv"
`include "wrGen.sv"
`include "rdGen.sv"
`include "interface.sv"
`include "wrBfm.sv"
`include "rdBfm.sv"
`include "wrMon.sv"
`include "rdMon.sv"
`include "wrCov.sv"
`include "rdCov.sv"
`include "wrAgent.sv"
`include "rdAgent.sv"
`include "sbd.sv"
`include "env.sv"
